module sr_latch(S,R,Q,Qbar);
input S,R;
output Q,Qbar;
nor N1(Q,S,Qbar);
nor N2(Qbar,R,Q);
endmodule