module encoder_8to3(A7,A6,A5,A4,A3,A2,A1,A0,B,C,D);
input A7,A6,A5,A4,A3,A2,A1,A0;
output B,C,D;

assign B=(A4|A5|A6|A7);
assign C=(A2|A3|A6|A7);
assign D=(A1|A3|A5|A7);

endmodule