module mux_16to1(in,sel,out);
input [15:0]in;
input[0:3]sel;
output out;
assign out=in[sel];
endmodule